library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity RippleCPU is
end RippleCPU;

architecture Behavioral of RippleCPU is

begin


end Behavioral;
